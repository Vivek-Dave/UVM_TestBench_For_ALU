
interface intf();
    // ------------------- port declaration-------------------------------------
    logic [7:0] in1;
    logic [7:0] in2;
    logic [3:0] s;
    logic m;
    logic cin;

    logic [7:0] out;
    logic cout;
    logic aeb;
    //--------------------------------------------------------------------------
    //--------------------------------------------------------------------------
        
endinterface

