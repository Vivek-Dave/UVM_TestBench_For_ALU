
`include "interface.sv"
`include "tb_pkg.sv"
module top;
  import uvm_pkg::*;
  import tb_pkg::*;
  
  //----------------------------------------------------------------------------
  intf i_intf();
  //----------------------------------------------------------------------------

  //----------------------------------------------------------------------------
  alu DUT(.in1 (i_intf.in1),
          .in2 (i_intf.in2),
          .s   (i_intf.s),
          .m   (i_intf.m),
          .cin (i_intf.cin),
          .out (i_intf.out),
          .cout(i_intf.cout),
          .aeb (i_intf.aeb)
          );
  //----------------------------------------------------------------------------               
  
  //----------------------------------------------------------------------------
  initial begin
    $dumpfile("dumpfile.vcd");
    $dumpvars;
  end
  //----------------------------------------------------------------------------

  //----------------------------------------------------------------------------
  initial begin
    uvm_config_db#(virtual intf)::set(uvm_root::get(),"","vif",i_intf);
  end
  //----------------------------------------------------------------------------

  //----------------------------------------------------------------------------
  initial begin
    run_test("alu_test");
  end
  //----------------------------------------------------------------------------
endmodule

